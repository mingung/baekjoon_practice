module relu(convol, reluValue);
input convol;
output reluValue;

if (convol <= 0)
assign 
else
assign 
endmodule